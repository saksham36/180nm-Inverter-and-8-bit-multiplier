library verilog;
use verilog.vl_types.all;
entity multiply_tb is
end multiply_tb;
